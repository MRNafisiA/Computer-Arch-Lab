module instruction_memory(address, instruction);
    input [41:0] address;
    output [31:0] instruction;

//      instrudction must be set here!
//    assign instruction = ;

endmodule